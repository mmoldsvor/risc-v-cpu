package cpu_package;
    typedef enum {
        ADD = 3'b000,
        SUB = 3'b001,
        AND = 3'b010,
        OR  = 3'b011
    } alu_function_t;
endpackage